dshultz@SURF.37